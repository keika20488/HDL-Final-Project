// map
module draw_map(
    input [3:0] state,
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    input isLocked,
    output reg [16:0] pixel_addr,
    output reg isObject
);
parameter [3:0] STAGE1 = 2, STAGE2 = 4, STAGE3 = 6;

parameter [0:40] map [0:40] = {
    41'b11111111111111111111111111111111111111111,
    41'b10000000000000000000000000000000000000001,
    41'b10000000000000000000000000000000000000001,
    41'b10000000000000000000000000000000000000001,
    41'b10001111111111111110001111111111111110001,
    41'b10001111111111111110001111111111111110001,
    41'b10001111111111111110001111111111111110001,
    41'b10001110000000000000000000000000001110001,
    41'b10001110000000000000000000000000001110001,
    41'b10001110000000000000000000000000001110001,
    41'b10001110001111111111111111111110001110001,
    41'b10001110001111111111111111111110001110001,
    41'b10001110001111111111111111111110001110001,
    41'b10001110000000000000000000000000001110001,
    41'b10001110000000000000000000000000001110001,
    41'b10001110000000000000000000000000001110001,
    41'b10001110001111111111111111111111111110001,
    41'b10001110001111111111111111111111111110001,
    41'b10001110001111111111111111111111111110001,
    41'b10001110000000000000000000000000000000000,
    41'b10001110000000000000000000000000000000000,
    41'b10001110000000000000000000000000000000000,
    41'b10001110001111111111111111111111111110001,
    41'b10001110001111111111111111111111111110001,
    41'b10001110001111111111111111111111111110001,
    41'b10001110001110000000000000000000001110001,
    41'b10001110001110000000000000000000001110001,
    41'b10001110001110000000000000000000001110001,
    41'b10001110001110001110001110001110001110001,
    41'b10001110001110001110001110001110001110001,
    41'b10001110001110001110001110001110001110001,
    41'b10000000000000001110001110001110001110001,
    41'b10000000000000001110001110001110001110001,
    41'b10000000000000001110001110001110001110001,
    41'b11111111111111111111111110001110001110001,
    41'b11111111111111111111111110001110001110001,
    41'b11111111111111111111111110001110001110001,
    41'b10000000000000000000000000001110000000001,
    41'b10000000000000000000000000001110000000001,
    41'b10000000000000000000000000001110000000001,
    41'b11111111111111111111111111111111111111111
};
//41=1+39+1
//205*205
wire [8:0] x,y;
assign x = h_cnt>>1;
assign y = v_cnt>>1;
always@(*)begin
    isObject = 0;
    pixel_addr = 0;
    case(state)
    STAGE1, STAGE2, STAGE3:begin
        if(x >= 260 && x <270 && y>=127 && y<137)begin
            if(isLocked)begin
                pixel_addr = (x + 80 + (y - 107)*360)%86400;
                isObject = 1;
            end else begin
                pixel_addr = (x + 90 + (y - 107)*360)%86400;
                isObject = 1;
            end
        end else if(x >= 60 && x < 265 && y >= 30 && y < 235)begin
            if(map[(y - 30)/5][(x - 60)/5])begin
                pixel_addr = (x%5 + 330 + (y%5 + 30) * 360)%86400;
                isObject = 1;
            end 
        end
    end
    endcase
end
endmodule