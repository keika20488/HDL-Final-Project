// wall
module draw_map(
    input [3:0] state,
    input [9:0] h_cnt,
    input [9:0] v_cnt,
    output reg [16:0] pixel_addr,
    output reg isObject
);
parameter [3:0] TITLE = 0, STAFF = 1;
parameter [3:0] STAGE1 = 2, SUCCESS1 = 3;
parameter [3:0] STAGE2 = 4, SUCCESS2 = 5;
parameter [3:0] STAGE3 = 6, SUCCESS3 = 7, FAIL = 8;

parameter [0:40] map [0:40] = {
41'b11111111111111111111111111111111111111111,
41'b10000000000000000000000000000000000000001,
41'b10000000000000000000000000000000000000001,
41'b10000000000000000000000000000000000000001,
41'b10001111111111111110001111111111111110001,
41'b10001111111111111110001111111111111110001,
41'b10001111111111111110001111111111111110001,
41'b10001110000000000000000000000000001110001,
41'b10001110000000000000000000000000001110001,
41'b10001110000000000000000000000000001110001,
41'b10001110001111111111111111111110001110001,
41'b10001110001111111111111111111110001110001,
41'b10001110001111111111111111111110001110001,
41'b10001110000000000000000000000000001110001,
41'b10001110000000000000000000000000001110001,
41'b10001110000000000000000000000000001110001,
41'b10001110001111111111111111111111111110001,
41'b10001110001111111111111111111111111110001,
41'b10001110001111111111111111111111111110001,
41'b10001110000000000000000000000000000000000,
41'b10001110000000000000000000000000000000000,
41'b10001110000000000000000000000000000000000,
41'b10001110001111111111111111111111111110001,
41'b10001110001111111111111111111111111110001,
41'b10001110001111111111111111111111111110001,
41'b10001110001110000000000000000000001110001,
41'b10001110001110000000000000000000001110001,
41'b10001110001110000000000000000000001110001,
41'b10001110001110001110001110001110001110001,
41'b10001110001110001110001110001110001110001,
41'b10001110001110001110001110001110001110001,
41'b10000000000000001110001110001110001110001,
41'b10000000000000001110001110001110001110001,
41'b10000000000000001110001110001110001110001,
41'b11111111111111111111111110001110001110001,
41'b11111111111111111111111110001110001110001,
41'b11111111111111111111111110001110001110001,
41'b10000000000000000000000000001110000000001,
41'b10000000000000000000000000001110000000001,
41'b10000000000000000000000000001110000000001,
41'b11111111111111111111111111111111111111111
};
//41=1+39+1
//205*205
wire [8:0] x,y;
assign x = h_cnt>>1;
assign y = v_cnt>>1;
always@(*)begin
    isObject = 0;
    pixel_addr = 0;
    case(state)
    STAGE1, STAGE2, STAGE3:begin
        if(x >= 60 && x < 265 && y >= 30 && y < 235)begin
            if(map[(y - 30)/5][(x - 60)/5])begin
                pixel_addr = (x%5 + 330 + (y%5 + 30) * 360)%86400;
                isObject = 1;
            end 
        end
    end
    endcase
    
end
endmodule
//200*200->40*40 player20*20->4*4
/*

111111111111111111111111111111111111111
100000000000000000010000000000000000001
100000000000000000010000000000000000001
100000000000000000010000000000000000001
100000000000000000010000000000000000001
100001111111111000011111111111111100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000011111111111111111110000100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000011111111111111111111111100001
100001000000000000000000000000000000000
100001000000000000000000000000000000000
000001000000000000000000000000000000000
000001000000000000000000000000000000000
000001000011111111111111111111111100001
000001000010000000000000000000000100001
100001000010000000000000000000000100001
100001000010000000000000000000000100001
100001000010000000000000000000000100001
100001000010000100001100001000000100001
100001000010000100001100001000000000001
100001000010000100001100001000000000001
100001000010000100001100001000000000001
100000000000000100001100001000000000001
100000000000000100001100001000011100001
100000000000000100001100001000011100001
100000000000000100001100001000011100001
111111111111111111111100001000011100001
111111111111111111111100001000011100001
100000000000000000000000001000000000001
100000000000000000000000001000000000001
100000000000000000000000001000000000001
100000000000000000000000001000000000001
111111111111111111111111111111111111111

11111111111111111111111111111111111111111
10000000000000000000000000000000000000001
10000000000000000000000000000000000000001
10000000000000000000000000000000000000001
10001111111111111000001111111111111000001
10001000000000000000000000000000001000001
10001000000000000000000000000000001000001
10001000000000000000000000000000001000001
10001000000000000000000000000000001000001
10001000000000000000000000000000001000001
10001000001111111111111111111000001000001
10001000000000000000000000000000001000001
10001000000000000000000000000000001000001
10001000000000000000000000000000001000001
10001000000000000000000000000000001000001
10001000000000000000000000000000001000001
10001000001111111111111111111111111000001
10001000000000000000000000000000000000001
10001000000000000000000000000000000000001
10001000000000000000000000000000000000001
10001000000000000000000000000000000000001
10001000000000000000000000000000000000001
10001000001111111111111111111111111000001
10001000001000000000000000000000001000001
10001000001000000000000000000000001000001
10001000001000000000000000000000001000001
10001000001000000000000000000000001000001
10001000001000000000000000000000001000001
10001000001000001000001000001000001000001
10000000000000001000001000001000001000001
10000000000000001000001000001000001000001
10000000000000001000001000001000001000001
10000000000000001000001000001000001000001
10000000000000001000001000001000001000001
11111111111111111111111000001000001000001
10000000000000000000000000001000000000001
10000000000000000000000000001000000000001
10000000000000000000000000001000000000001
10000000000000000000000000001000000000001
10000000000000000000000000001000000000001
11111111111111111111111111111111111111111
*/