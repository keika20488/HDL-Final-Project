`define rec_h = 20;
`define rec_v = 20;
module game_play (
    input rst,
    input clk,
    inout wire PS2_DATA,
    inout wire PS2_CLK,
    output reg [1:0] todo,
    output reg [3:0] state,
    output reg [3:0] player_state,
    output reg [3:0] boss_state,
    output reg [8:0] player_x,
    output reg [8:0] player_y,
    output reg [8:0] boss_x,
    output reg [8:0] boss_y,
    output reg [8:0] obj_x,
    output reg [8:0] obj_y,
    output reg [1:0] key_find,
    output reg [3:0] play_valid,
    output reg isDark
);

// Keyboard
wire [130:0] key_down;
wire [6:0] last_change;
reg [4:0] key_num;

KeyboardDecoder key_de (
    .key_down(key_down),
    .last_change(last_change),
    .key_valid(been_ready),
    .PS2_DATA(PS2_DATA),
    .PS2_CLK(PS2_CLK),
    .rst(rst),
    .clk(clk)
);

// KeyCodes: n, b, r, 1-3, WASD, right shift
parameter [6:0] KEY_CODES [0:10] = {
    7'b101_1001,  //right shift//59
    7'b110_1001,  //1          //69
    7'b111_0010,  //2          //72
    7'b111_1010,  //3          //7A
    7'b001_1101,  //w  //up    //1D
    7'b001_1100,  //a  //left  //1C
    7'b001_1011,  //s  //down  //1B
    7'b010_0011,  //d  //right //23
    7'b011_0001,  //n  //next  //31
    7'b011_0010,  //b  //back  //32
    7'b010_1101   //r  //retry //2D
};

always @(*) begin
    case(last_change)
    KEY_CODES[0] : key_num = 0;
    KEY_CODES[1] : key_num = 1;
    KEY_CODES[2] : key_num = 2;
    KEY_CODES[3] : key_num = 3;
    KEY_CODES[4] : key_num = 4;
    KEY_CODES[5] : key_num = 5;
    KEY_CODES[6] : key_num = 6;
    KEY_CODES[7] : key_num = 7;
    KEY_CODES[8] : key_num = 8;
    KEY_CODES[9] : key_num = 9;
    KEY_CODES[10]: key_num = 10;
    default : key_num = 15;
    endcase
end


// State: title, stage1, success1, stage2, success2, stage3, success3, fail3, staff
parameter [3:0] TITLE = 0, STAFF = 1;
parameter [3:0] STAGE1 = 2, SUCCESS1 = 3;
parameter [3:0] STAGE2 = 4, SUCCESS2 = 5;
parameter [3:0] STAGE3 = 6, SUCCESS3 = 7, FAIL = 8;
reg pass, fail;

always @(posedge clk or posedge rst) begin
    if (rst) play_valid <= 4'b0010;
    else begin
        case(state)
        SUCCESS1: play_valid <= 4'b0110;
        SUCCESS2: play_valid <= 4'b1110;
        default: play_valid <= 4'b1111;
        endcase
    end
end

always @(posedge clk or posedge rst) begin
    if (rst) state <= TITLE;
    else begin
        case(state)
        TITLE: begin
            if (key_down[last_change] && key_num < 4 && play_valid[key_num])
                state <= key_num * 2;
            else state <= TITLE;
        end
        STAGE1: begin
            if (pass) state <= SUCCESS1;
            else state <= STAGE1;
        end
        SUCCESS1: begin
            if (key_down[last_change]) begin
                if (key_num == 8) state <= STAGE2;
                else if (key_num == 9) state <= TITLE;
                else state <= SUCCESS1;
            end else state <= SUCCESS1;
        end
        STAGE2: begin
            if (pass) state <= SUCCESS2;
            else state <= STAGE2;
        end
        SUCCESS2: begin
            if (key_down[last_change]) begin
                if (key_num == 8) state <= STAGE3;
                else if (key_num == 9) state <= TITLE;
                else state <= SUCCESS2;
            end else state <= SUCCESS2;
        end
        STAGE3: begin
            if (pass) state <= SUCCESS3;
            else if (fail) state <= FAIL;
            else state <= STAGE3;
        end
        SUCCESS3: begin
            if (key_down[last_change] && key_num == 8)
                state <= STAFF;
            else state <= SUCCESS3;
        end
        FAIL: begin
            if (key_down[last_change]) begin
                if (key_num == 10) state <= STAGE3;
                else if (key_num == 9) state <= TITLE;
                else state <= FAIL;
            end else state <= FAIL;
        end
        STAFF: begin
            if (key_down[last_change] && key_num == 9)
                state <= TITLE;
            else state <= STAFF;
        end
        default: state <= state;
        endcase
    end
end

// Todo: key, light, door
parameter [1:0] NONE = 0, FIND_KEY = 1, FIND_LIGHT = 2, FIND_DOOR = 3;

always @(posedge clk or posedge rst) begin
    if (rst) todo <= NONE;
    else begin
        case(state)
        STAGE1: begin
            if (key_find < 3) todo <= FIND_KEY;
            else todo <= FIND_DOOR;
        end
        STAGE2: begin
            if (isDark) todo <= FIND_LIGHT;
            else if (key_find < 3) todo <= FIND_KEY;
            else todo <= FIND_DOOR;
        end
        STAGE3: begin
            if (key_find < 3) todo <= FIND_KEY;
            else todo <= FIND_DOOR;
        end
        default: todo <= NONE;
        endcase
    end
end


// Clock Divider
clock_divider #(23) div_23(.clk(clk), .clk_div(clk_23));

// Player Position
parameter [3:0] UP1 = 0, UP2 = 1, UP3 = 2;
parameter [3:0] RIGHT1 = 3, RIGHT2 = 4, RIGHT3 = 5;
parameter [3:0] LEFT1 = 6, LEFT2 = 7, LEFT3 = 8;
parameter [3:0] DOWN1 = 9, DOWN2 = 10, DOWN3 = 11;

parameter [40:0] map [0:40] = {
41'b11111111111111111111111111111111111111111,
41'b10000000000000000000000000000000000000001,
41'b10000000000000000000000000000000000000001,
41'b10000000000000000000000000000000000000001,
41'b10001111111111111000001111111111111000001,
41'b10001000000000000000000000000000001000001,
41'b10001000000000000000000000000000001000001,
41'b10001000000000000000000000000000001000001,
41'b10001000000000000000000000000000001000001,
41'b10001000000000000000000000000000001000001,
41'b10001000001111111111111111111000001000001,
41'b10001000000000000000000000000000001000001,
41'b10001000000000000000000000000000001000001,
41'b10001000000000000000000000000000001000001,
41'b10001000000000000000000000000000001000001,
41'b10001000000000000000000000000000001000001,
41'b10001000001111111111111111111111111000001,
41'b00001000000000000000000000000000000000001,
41'b00001000000000000000000000000000000000001,
41'b00001000000000000000000000000000000000001,
41'b00001000000000000000000000000000000000001,
41'b00001000000000000000000000000000000000001,
41'b10001000001111111111111111111111111000001,
41'b10001000001000000000000000000000001000001,
41'b10001000001000000000000000000000001000001,
41'b10001000001000000000000000000000001000001,
41'b10001000001000000000000000000000001000001,
41'b10001000001000000000000000000000001000001,
41'b10001000001000001000001000001000001000001,
41'b10000000000000001000001000001000001000001,
41'b10000000000000001000001000001000001000001,
41'b10000000000000001000001000001000001000001,
41'b10000000000000001000001000001000001000001,
41'b10000000000000001000001000001000001000001,
41'b11111111111111111111111000001000001000001,
41'b10000000000000000000000000001000000000001,
41'b10000000000000000000000000001000000000001,
41'b10000000000000000000000000001000000000001,
41'b10000000000000000000000000001000000000001,
41'b10000000000000000000000000001000000000001,
41'b11111111111111111111111111111111111111111
};

always @(posedge clk_23 or posedge rst) begin
    if (rst) player_state <= RIGHT1;
    else begin
        case(state)
        STAGE1, STAGE2, STAGE3: begin
            if(key_down[last_change]) begin
                case (key_num)
                4: player_state <= (player_state == UP2) ? UP3 : UP2;
                5: player_state <= (player_state == LEFT2) ? LEFT3 : LEFT2;
                6: player_state <= (player_state == DOWN2) ? DOWN3 : DOWN2;
                7: player_state <= (player_state == RIGHT2) ? RIGHT3 : RIGHT2;
                default: player_state <= player_state;
                endcase
            end else player_state <= player_state / 3 * 3;
        end
        default: player_state <= RIGHT1;
        endcase
    end
end

always @(posedge clk_23) begin
    player_x <= player_x;
    player_y <= player_y;
    case(state)
    STAGE1, STAGE2, STAGE3: begin
        if(key_down[last_change]) begin
            case (key_num)
            4: begin
                if(!map[(player_y -1 - 30)/5][(player_x - 60)/5] && !map[(player_y -1 - 30 +10)/5][(player_x - 60 +10)/5])begin
                    player_y <= player_y - 1;
                end
            end
            5: begin
                if(!map[(player_y - 30)/5][(player_x -1 - 60)/5] && !map[(player_y - 30 +10)/5][(player_x -1 - 60 +10)/5])begin
                    player_x <= player_x - 1;
                end
            end
            6: begin
                if(!map[(player_y +1 - 30)/5][(player_x - 60)/5] && !map[(player_y +1 - 30 +10)/5][(player_x - 60 +10)/5])begin
                    player_y <= player_y + 1;
                end
            end
            7: begin
                if(!map[(player_y - 30)/5][(player_x +1 - 60)/5] && !map[(player_y - 30 +10)/5][(player_x +1 - 60 +10)/5])begin
                    player_x <= player_x + 1;
                end
            end
            endcase
        end
    end
    default: begin
        player_x <= 65;
        player_y <= 125;
    end
    endcase
end
//Boss position
reg [8:0] next_boss_x;
reg [8:0] next_boss_y;

parameter [337:0] shortest_dir[0:168]={
338'b00101010101010101010101010010000000000100000000000100100101010101010101010001001001000000000000000100010010010101010101010101000100100100000000000000000001001001010101010101010101010010001000000000000000000100100010001010101010101001001000100010001000100010010010101010100010001000100100000000000000000010001001001010101010101010100101010,
338'b11001010101010101010101010111111111111101111111111101111101010101010101010111011111011111111111111101110111110101010101010101011101111101111111111111111111011111010101010101010101010111110111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111110111011111111111111111111101010,
338'b11110010101010101010101010111111111111101111111111101111101010101010101010111011111011111111111111101110111110101010101010101011101111101111111111111111111011111010101010101010101010111110111111111111111111101111101111111111111111111011111111111111111111111110111111111111111111111011101111111111111111111110111011111111111111111111101010,
338'b11111100101010101010101010111111111111101111111111101111101010101010101010111011111011111111111111101110111110101010101010101011101111101111111111111111111011111010101010101010101010111110111111111111111111101111101111111111111111111011111011111111111111101110111111111111111111111011101111111111111111111110111011111111111111111111101010,
338'b11111111001010101010101010111111111111101111111111101111101010101010101010111011111011111111111111101110111110101010101010101011101111101111111111111111111011111010101010101010101010111110111111111111111111101111101110101010101010111011111011101110111011101110111110101011101110111011101111111111111111101110111010101010101010101011101010,
338'b11111111110010101010101010111111111111101111111111101111101010101010101010111011111011111111111111101110111110101010101010101011101111101111111111111111111011111010101010101010101010111110111111111111111111101111101110101010101010111011111011101110111011101110111010101011101110111011101111111111111111101110111010101010101010101011101010,
338'b11111111111100101010101010111111111111011111111111101111010101010101010101111011110111111111111111011110111101010101010101010111101111011111111111111111111011110101010101011010101010111101111111111111111111101111011101010101010110111011110111011101110111101110010101010111011101111011101111111111111111011110111001010101010101010111101010,
338'b11111111111111001010101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111111101010101010111111111111111111111111101111111111111111111010111011111111111111111111101110111111111111111111111011101111111111111111111110111011111111111111111111101010,
338'b11111111111111110010101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111110101010101010111111111111111111111111101111111111111111101010111011111111111111111011101110111111111111111110111011101111111111111111101110111010101010101010101011101010,
338'b11111111111111111100101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111010101010101010111111111111111111111111101111111111111110101010111011111111111111111011101110111111111111111110111011101111111111111111101110111010101010101010101011101010,
338'b11111111111111111111001010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111101010101010101010111111111111111111111111101111111111111010101010111011111111111110111011101110111111111111101110111011101111111111111111101110111010101010101010101011101010,
338'b11111111111111111111110010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111110101010101010101010111111111111111111111111101111111111101010101010111011111111111110111011101110111111111111101110111011101111111111111111101110111010101010101010101011101010,
338'b11111111111111111111111100111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111111111111111110111110101010101010101010101111101111111111111111111011111011101010101010101110111110111011101110111011101010101010111011101110111011111111111111111011101110101010101010101010111010101,
338'b00000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000010000000000000000000000000100000000000000000000000001000101010101010100000000010001000000000000000000000100010001010101010101000001000100010001000100010000010101010100010001000100000000000000000000010001000001010101010101010100010000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000010101010101010101000000000100000000000000010000000001010101010101010100000000010000000000000000000000000101010101010100000000000001000000000000000000000000010001010101010101000000000100010001000100000000010101010100010001000000000000000000000000010000000001010101010101010100000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001000000000000000000000000010000000000000000000000000100000101010101010101010101000001000000000000000000010000010001010101010101000100000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000000000000000000000100010000000000000000000001000101010101010101000000010001000000000000000000000100010001010101010101000001000100010001000100010000010101010100010001000100000000000000000000010001000001010101010101010100010100,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b10101010101010101010101010101010101010101010101010101010001010101010101010101010100110101010101010101010101001010101010101011010100110011010101010101010100101100101010101010101010101011001101010101010101010010110011001010101010101100101100110011001100110011001010101010110011001100110011010101010101010011001100101010101010101010110010101,
338'b10101010101010101010101010101010101010101010101010101010110010101010101010101010101110101010101010101010101011111111111111101010101010111010101010101010101011101111111111111111111111111011101010101010101010111110111011111111111111101111101110111011101110111011111111111110111011101110111010101010101010111011101111111111111111111110111111,
338'b10101010101010101010101010101010101010101010101010101010111100101010101010101010101110101010101010101010101011111111111110101010101010111010101010101010101010101111111111111111111110111011101010101010101010101110111011111111111111101011101110111011101110111010111111111110111011101110101010101010101010111011101011111111111111111110101010,
338'b10101010101010101010101010101010101010101010101010101010111111001010101010101010101110101010101010101010101011111111111010101010101010111010101010101010101010101111111111111111111010101011101010101010101010101110111011111111111111101011101110111011101110111010111111111110111011101110101010101010101010111010101011111111111111111110101010,
338'b00000000000000000000000000000000000000000000000000000000111111110010101010000000001100000000000000100000000011111111101010101000000000110000000000000000000000001111111111111111000000000011000000000000000000000000110011111111111111000011001100110011001100110000111111111100110011000000000000000000000000110000000011111111111111111100000000,
338'b11111111111111111111111111111111111111111111111111111111111111111100101010111111111111111111111111101111111111111110101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
338'b11111111111111111111111111111111111111111111111111111111111111111111001010111111111111111111111111101111111111111010101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
338'b11111111111111111111111111111111111111111111111111111111111111111111110010111111111111111111111111101111111111101010101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
338'b11111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111011111111101010101010101010111111111011111111111111111111111110101010101010101011111111101111111111111111111110111011101010101010101111101110111011101110111011111010101010111011101110111111111111111111111011111111101010101010101010111111111,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000010000000000000000000100000101010101010101010101000001000000000000000000010000010001010101010101000101000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001010101010000000000000100010000000000000000000001000101010101010101010000010001000000000000000000000100010001010101010101000001000100010001000100010000010101010100010001000100000000000000000000010001000001010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001010101010101010100010100010000000000000000000101000101010101010101010101010001000000000000000000010100010001010101010101000101000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010100000000010000000000000000000000000101010101010101010000000001000000000000000000000100010001010101010101000001000100010001000100010000010101010100010001000100000000000000000000010000000001010101010101010100000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010000000000010000010000000000000000000100000101010101010101010101000001000000000000000000010100010001010101010101000101000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001010101010100000000000100010000000000000000000001000101010101010101010100010001000000000000000000000100010001010101010101000001000100010001000100010000010101010100010001000100000000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000100001010000101010101010101000010100010000000000000000000101000101010101010101010101010001000000000000000000010100010001010101010101000101000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b11111111111111111111111111111111111111111111111111111111111111111111111010111111111111111111111111101111111111001010101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
338'b11111111111111111111111111111111111111111111111111111111111111111111101010111111111111111111111111101111111111110010101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
338'b11111111111111111111111111111111111111111111111111111111111111111110101010111111111111111111111111101111111111111100101010101011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
338'b10101010101010101010101010101010101010101010101010101010111111111010101010101011101110101010101010101011111011111111001010101010111110111010101010101010101111101111111111111111111111111011101010101010101010111110111011111111111111101111101110111011101110111011111111111110111011101110111010101010101010111011101111111111111111111110111111,
338'b10101010101010101010101010101010101010101010101010101010111111101010101010101010101110101010101010101010111011111111110010101010111110111010101010101010101111101111111111111111111111111011101010101010101010111110111011111111111111101111101110111011101110111011111111111110111011101110111010101010101010111011101111111111111111111110111111,
338'b10101010101010101010101010101010101010101010101010101010111110101010101010101010101110101010101010101010101011111111111100101010101110111010101010101010101111101111111111111111111111111011101010101010101010111110111011111111111111101111101110111011101110111011111111111110111011101110111010101010101010111011101111111111111111111110111111,
338'b10101010101010101010101010101010101010101010101010101010111010101010101010101010101110101010101010101010101011111111111111001010101010111010101010101010101011101111111111111111111111111011101010101010101010111110111011111111111111101111101110111011101110111011111111111110111011101110111010101010101010111011101111111111111111111110111111,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000011111111111111110000000000110000000000000000000000001111111111111111111100110011000000000000000000001100110011111111111111000011001100110011001100110000111111111100110011001100000000000000000000110011000011111111111111111100000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000001010101010100000000000000010000000000000000000100000101010101010101010101010001000000000000000000010100010001010101010101000101000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000001010101010101000000000000010000000000000000000001000101010101010101010101010001000000000000000000010100010001010101010101000101000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000100000000000000000000000101000000000000000000000001010000000000000000000000010100000000000000000000000101000101010101010101010101010001000000000000000000010100010001010101010101000101000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000001010101010101000000000000010000000000000000000001000101010101010101010101010001000000000000000000010100010001010101010101000101000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000010100000000000000000000000100000000000000000000000001010101010101010000000000010000000000000000000100000101010101010101010101010001000000000000000000010100010001010101010101000101000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000010000000000000000000000100100000000000000000000001001000000000000000000000010010000000000000000000000100100000000000000000000001001000010101010101010101010010001000000000000000000100100010001010101010101001001000100010001000100010010010101010100010001000100100000000000000000010001001001010101010101010100101010,
338'b11111111111111111111111010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111100101010101010101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111110111011111111111111111111101010,
338'b11111111111111111111101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111001010101010101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111011101111111111111111111110111011111111111111111111101010,
338'b11111111111111111110101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111110010101010101010111111111111111111111111101111111111111111111111111011111111111111111111101110111111111111111111111011101111111111111111111110111011111111111111111111101010,
338'b11111111111111111010101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111100101010101010111111111111111111111111101111111111111111111110111011111111111111111111101110111111111111111111111011101111111111111111111110111011111111111111111111101010,
338'b11111111111111101010101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111111001010101010111111111111111111111111101111111111111111111010111011111111111111111111101110111111111111111111111011101111111111111111111110111011111111111111111111101010,
338'b10101010101010101010101010111010101010111010101010101110111111111111111111101011101110101010101010111010111011111111111111111110101110111010101010101010101011101111111111110010101010111011101010101010101010101110111011111111101010101011101110111011101010101010111111111110111010101010101010101010101010101010101010101010101010101010101010,
338'b10101010101010101010101010101010101010101010101010101110111111111111111111101011101110101010101010111010111011111111111111111110101110111010101010101010101011101111111111111100101010111011101010101010101010101110111011111110101010101011101110111011101010101010111111111110111010101010101010101010101010101010101010101010101010101010101010,
338'b10101010101010101010101010101010101010101010101010101010111111111010101010101011101110101010101010111010111011111111111111111110101110111010101010101010101011101111111111111111001010111011101010101010101010101110111011111010101010101011101110111010101010101010111111111110101010101010101010101010101010101010101010101010101010101010101010,
338'b10101010101010101010101010101010101010101010101010101010111111101010101010101010101110101010101010101010111011111111111111111110101110111010101010101010101011101111111111111111110010111011101010101010101010101110111011101010101010101011101110111010101010101010111111111110101010101010101010101010101010101010101010101010101010101010101010,
338'b00000000000000000000000000000000000000000000000000000000111100000000000000000000001100000000000000000000000011111111111111110000001100110000000000000000000011001111111111111111111100110011000000000000000000011100110001010101010101000111001100110001000100010001111111111100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000010101000000000000000000000100000000000000000000000001010101010101010100010000010000000000000000000100000101010101010101010101000001000000000000000000010100010001010101010101000101000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b01000000000000000000000000010101010101000101010101000101000000000000000000010001010001010101010101000100010100000000000000000001000101000101010101010101010001010000000000000000000000010100010101010101010101000101010101010101010101010001010101010101010101010100010101010101010101010101000101010101010101010101010001010101010101010101010000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101000100000000000001000100010001000000000000010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000010101010000000000000000000100000000000000010001000001010101010101010100010000010000000000000000000100000101010101010101010101000001000000000000000000010000010001010101010101000101000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b01010000000000000000000000010101010101000101010101000101000000000000000000010001010001010101010101000100010100000000000000000001000101000101010101010101010001010000000000000000000000010100010101010101010101000101000101010101010101010001010101010101010101010100010101010101010101010101000101010101010101010101010001010101010101010101010100,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b01010101010101010101010110010101010101010101010101100101010101010101010101011001010101010101010101010110010101010101010101010101100101010101010101010101011001010101010101010101010110010101010101010101010101100101010100101010101010011001010101010110011001100110010101010101100110011001100101010101010101100110011010101010101010101001101010,
338'b11111111111111111111111010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111111111111111010111111111111111111111111101111111111001010101010111011111111111110111011101110111111111111101110111011101111111111111111101110111010101010101010101011101010,
338'b11111111111111111111101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111111111111101010111111111111111111111111101111111111110010101010111011111111111101111011101110111111111111011110111011101111111111111111101110111010101010101010101011101010,
338'b11111111111111111110101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111111111110101010111111111111111111111111101111111111111100101010111011111111111111111011101110111111111111111110111011101111111111111111101110111010101010101010101011101010,
338'b11111111111111111010101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111111111010101010111111111111111111111111101111111111111111001010111011111111111111110111101110111111111111111101111011101111111111111111011110111001010101010101010111101010,
338'b11111111111111101010101010111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111111101010101010111111111111111111111111101111111111111111110010111011111111111111111111101110111111111111111111111011101111111111111111111110111011111111111111111111101010,
338'b11111111010101010101010101111111111111111111111111011111111111111111111111110111111111111111111111111101111111111111111111111111011111111111111111111111110111111111111101010101010101111111111111111111111111011111111111111111111100110111111111111111111111011101111111111111111111110111011111111111111111111101110111111111111111111111010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101000000000000010001000100010001000000000000010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000010101010101010101000100000100000000000000010001000001010101010101010100010000010000000000000000000100000101010101010101010101000001000000000000000000010000010001010101010101000100000100010001000100010001010101010100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b01010100000000000000000000010101010101000101010101000101000000000000000000010001010001010101010101000100010100000000000000000001000101000101010101010101010001010000000000000000000000010100010101010101010101000101000101010101010101010001010001010101010101010100010101010101010101010101000101010101010101010101010001010101010101010101010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b01010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010100000000000000010001010101000100010001000100010101010101000100010001000101010101010101000100010000000000000000000001000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010000000001010101010101010100000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000010101010101010101000000000000000000000000010000000000000000000000000100000000000000000000000001000000000000000000000000010000000000000000000000000100000000000001010101010101000000000000000000000000010000000000000000000000000100000000000000000000000001000000000000000000000100010000000000000000000001000100000000000000000000010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101000000000000010001000100010000000000000100010001000100010000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000100000000000100000101010101010101010001000001000000000000000100010000010101010101010101000100000100000000000000000001000001010101010101010101010000010000000000000000000100000100010101010101010001000001000100010001000100010001010101000100010001000100000000000000000100010001010101010101010101000101010,
338'b11111111111010101010101010111111111111101111111111101111101010101010101010111011111011111111111111101110111110101010101010101011101111101111111111111111111011111010101010101010101010111110111111111111111111101111101110101010101010111011111011101110111011101110110010101011101110111011101111111111111111101110111010101010101010101011101010,
338'b11111111000000000000000000111111111111001111111111001111000000000000000000110011110011111111111111001100111100000000000000000011001111001111111111111111110011110000000000000000000000111100111111111111111111001111001110101010101010110011110011101110111011101100111100101011101110111011001111111111111111101110111010101010101010101011101010,
338'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110101010101010111111111111101110111011101110111111001011101110111011101111111111111111101110111010101010101010101011101010,
338'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000110011111111001100110011001100111111110011001100110011001111111111111111001100110000000000000000000011000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001010101010101010100000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000001010101010101010101000000000000010000000000010000000000000000000000000100000000000000000000000001000000000000000000000000010000000000000000000000000100000000000101010101010101000000000000000000000000010000000000000000000000000100000000000000000000000001000000000000000000000000010000000000000000000001000100000000000000000000010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101000000000000010001000100010000000000010100010001000100000000000000000000010001000101010101010101010100010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010101010100000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000101010101010101010101000000000000010000000000010000000000000101010101000100000000000000000000000001000000000000000000000000010000000000000000000000000100000000010101010101010101000000000000000000000000010000000000000000000000000100000000000000000000000001000000000000000000000000010000000000000000000000000100000000000000000000010101,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101010100000000000000000000000000000000010101010000000000000000100000000000000000000000000001010101010101010000010101,
338'b10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000101010101010101010101010,
338'b10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011001010101010101010101010,
338'b10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011110010101010101010101010,
338'b10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011111100101010101010101010,
338'b10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011111111001010101010101010,
338'b10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011111111110010101010101010,
338'b10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011111111111100101010101010,
338'b10101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101011111111111111001010101010,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
338'b00101010101010101010101010000000000000100000000000100000000000101010101010001000000000000000000000100010000000000000000000000000100000000000000000000000001000000010101010101010101010000000000000000000000000100000000000000000000000001000000000000000000000000010000000000000000000000000100000000000000000000000001000000000000000000000001010,
338'b10101010101010101010101010101010101010101010101010101110101010101010101010101011101010101010101010101010111010101010101010101010101110101010101010101010101011101010101010101010101010111010101010101010101010101110111011111111111111101011101110111011101110111010111111111110111011101110101010101010101010111011101011111111111111111110110010,
338'b00000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000110000000000000000000000001100000000000000000000000011000000000000000000000000110000000000000000000000001100000011111111111111000011001100110011001100110000111111111100110011001100000000000000000000110011000011111111111111111100111100

};
wire [1:0] boss_dir;
assign boss_dir = {shortest_dir[(((player_x-60)/5)-1)/3*13+(((player_y-30)/5)-1)/3][((((boss_x-60)/5)-1)/3*13+(((boss_y-30)/5)-1)/3)*2+1],shortest_dir[(((player_x-60)/5)-1)/3*13+(((player_y-30)/5)-1)/3][((((boss_x-60)/5)-1)/3*13+(((boss_y-30)/5)-1)/3)*2]};

always @(posedge clk_23 or posedge rst) begin
    if (rst) boss_state <= RIGHT1;
    else begin
        case(state)
        STAGE3: begin
                case (boss_dir)
                0: boss_state <= (boss_state == UP2) ? UP3 : UP2;
                3: boss_state <= (boss_state == LEFT2) ? LEFT3 : LEFT2;
                1: boss_state <= (boss_state == DOWN2) ? DOWN3 : DOWN2;
                2: boss_state <= (boss_state == RIGHT2) ? RIGHT3 : RIGHT2;
                default: boss_state <= boss_state;
                endcase
        end
        default: boss_state <= RIGHT1;
        endcase
    end
end
always @(posedge clk_23 or posedge rst) begin
    if(rst)begin
        boss_x <=  250;
        boss_y <= 35;
    end
    else begin
        boss_x <=  250;
        boss_y <= 35;
        /*
        case(state)
        STAGE3:begin
        case(boss_dir)
            0:begin//up
                boss_x <= boss_x;
                boss_y <= boss_y - 1;
            end
            1:begin//down
                boss_x <= boss_x;
                boss_y <= boss_y + 1;
            end
            2:begin//right
                boss_x <= boss_x + 1;
                boss_y <= boss_y;
            end
            3:begin//left
                boss_x <= boss_x - 1;
                boss_y <= boss_y;
            end
            default:begin
                boss_x <= boss_x;
                boss_y <= boss_y;
            end
            endcase
            end
        endcase
        */
    end
end

// Object Position

// Collide
// Key
always @(posedge clk_23) begin
    key_find <= key_find;
    case(state)
    STAGE1, STAGE3: begin
        case (key_find)
        0: begin
            if (player_x >= 55 && player_x < 85 && player_y >= 25 && player_y < 55)
                key_find <= key_find + 1;
        end
        1: begin
            if (player_x >= 220 && player_x < 250 && player_y >= 25 && player_y < 55)
                key_find <= key_find + 1;
        end
        2: begin
            if (player_x >= 220 && player_x < 250 && player_y >= 195 && player_y < 255)
                key_find <= key_find + 1;
        end
        endcase
    end
    STAGE2: begin
        if (!isDark) begin
            case (key_find)
            0: begin
                if (player_x >= 55 && player_x < 85 && player_y >= 25 && player_y < 55)
                    key_find <= key_find + 1;
            end
            1: begin
                if (player_x >= 220 && player_x < 250 && player_y >= 25 && player_y < 55)
                    key_find <= key_find + 1;
            end
            2: begin
                if (player_x >= 220 && player_x < 250 && player_y >= 195 && player_y < 255)
                    key_find <= key_find + 1;
            end
            endcase
        end
    end
    default: key_find <= 0;
    endcase
end
// Pass
always @(posedge clk_23) begin
    if (key_find == 3 && player_x >= 250 && player_x < 280 && player_y >= 110 && player_y < 140)
        pass <= 1;
    else pass <= 0;
end
// Light
always @(posedge clk_23) begin
    isDark <= isDark;
    case(state)
    STAGE2: begin
        if (player_x >= 170 && player_x < 200 && player_y >= 125 && player_y < 150)
            isDark <= 0;
    end
    default: isDark <= 1;
    endcase
end
endmodule