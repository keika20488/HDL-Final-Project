`define rec_h = 20;
`define rec_v = 20;
module game_play (
    input rst,
    input clk,
    inout wire PS2_DATA,
    inout wire PS2_CLK,
    output reg [1:0] todo,
    output reg [3:0] state,
    output reg [3:0] player_state,
    output reg [3:0] boss_state,
    output reg [8:0] player_x,
    output reg [8:0] player_y,
    output reg [8:0] boss_x,
    output reg [8:0] boss_y,
    output reg [8:0] obj_x,
    output reg [8:0] obj_y,
    output reg [1:0] key_find,
    output reg [3:0] play_valid,
    output reg isDark
);

// Keyboard
wire [130:0] key_down;
wire [6:0] last_change;
reg [4:0] key_num;

KeyboardDecoder key_de (
    .key_down(key_down),
    .last_change(last_change),
    .key_valid(been_ready),
    .PS2_DATA(PS2_DATA),
    .PS2_CLK(PS2_CLK),
    .rst(rst),
    .clk(clk)
);

// KeyCodes: n, b, r, 1-3, WASD, right shift
parameter [6:0] KEY_CODES [0:10] = {
    7'b101_1001,  //right shift//59
    7'b110_1001,  //1          //69
    7'b111_0010,  //2          //72
    7'b111_1010,  //3          //7A
    7'b001_1101,  //w  //up    //1D
    7'b001_1100,  //a  //left  //1C
    7'b001_1011,  //s  //down  //1B
    7'b010_0011,  //d  //right //23
    7'b011_0001,  //n  //next  //31
    7'b011_0010,  //b  //back  //32
    7'b010_1101   //r  //retry //2D
};

always @(*) begin
    case(last_change)
    KEY_CODES[0] : key_num = 0;
    KEY_CODES[1] : key_num = 1;
    KEY_CODES[2] : key_num = 2;
    KEY_CODES[3] : key_num = 3;
    KEY_CODES[4] : key_num = 4;
    KEY_CODES[5] : key_num = 5;
    KEY_CODES[6] : key_num = 6;
    KEY_CODES[7] : key_num = 7;
    KEY_CODES[8] : key_num = 8;
    KEY_CODES[9] : key_num = 9;
    KEY_CODES[10]: key_num = 10;
    default : key_num = 15;
    endcase
end


// State: title, stage1, success1, stage2, success2, stage3, success3, fail3, staff
parameter [3:0] TITLE = 0, STAFF = 1;
parameter [3:0] STAGE1 = 2, SUCCESS1 = 3;
parameter [3:0] STAGE2 = 4, SUCCESS2 = 5;
parameter [3:0] STAGE3 = 6, SUCCESS3 = 7, FAIL = 8;
reg pass, fail;

always @(posedge clk or posedge rst) begin
    if (rst) play_valid <= 4'b0010;
    else begin
        case(state)
        SUCCESS1: play_valid <= 4'b0110;
        SUCCESS2: play_valid <= 4'b1110;
        default: play_valid <= play_valid;
        endcase
    end
end

always @(posedge clk or posedge rst) begin
    if (rst) state <= TITLE;
    else begin
        case(state)
        TITLE: begin
            if (key_down[last_change] && key_num < 4 && play_valid[key_num])
                state <= key_num * 2;
            else state <= TITLE;
        end
        STAGE1: begin
            if (pass) state <= SUCCESS1;
            else state <= STAGE1;
        end
        SUCCESS1: begin
            if (key_down[last_change]) begin
                if (key_num == 8) state <= STAGE2;
                else if (key_num == 9) state <= TITLE;
                else state <= SUCCESS1;
            end else state <= SUCCESS1;
        end
        STAGE2: begin
            if (pass) state <= SUCCESS2;
            else state <= STAGE2;
        end
        SUCCESS2: begin
            if (key_down[last_change]) begin
                if (key_num == 8) state <= STAGE3;
                else if (key_num == 9) state <= TITLE;
                else state <= SUCCESS2;
            end else state <= SUCCESS2;
        end
        STAGE3: begin
            if (pass) state <= SUCCESS3;
            else if (fail) state <= FAIL;
            else state <= STAGE3;
        end
        SUCCESS3: begin
            if (key_down[last_change] && key_num == 8)
                state <= STAFF;
            else state <= SUCCESS3;
        end
        FAIL: begin
            if (key_down[last_change]) begin
                if (key_num == 10) state <= STAGE3;
                else if (key_num == 9) state <= TITLE;
                else state <= FAIL;
            end else state <= FAIL;
        end
        STAFF: begin
            if (key_down[last_change] && key_num == 9)
                state <= TITLE;
            else state <= STAFF;
        end
        default: state <= state;
        endcase
    end
end

// Todo: key, light, door
parameter [1:0] NONE = 0, FIND_KEY = 1, FIND_LIGHT = 2, FIND_DOOR = 3;

always @(posedge clk or posedge rst) begin
    if (rst) todo <= NONE;
    else begin
        case(state)
        STAGE1: begin
            if (key_find < 3) todo <= FIND_KEY;
            else todo <= FIND_DOOR;
        end
        STAGE2: begin
            if (isDark) todo <= FIND_LIGHT;
            else if (key_find < 3) todo <= FIND_KEY;
            else todo <= FIND_DOOR;
        end
        STAGE3: begin
            if (key_find < 3) todo <= FIND_KEY;
            else todo <= FIND_DOOR;
        end
        default: todo <= NONE;
        endcase
    end
end


// Clock Divider
clock_divider #(23) div_23(.clk(clk), .clk_div(clk_23));

// Player Position
parameter [3:0] UP1 = 0, UP2 = 1, UP3 = 2;
parameter [3:0] RIGHT1 = 3, RIGHT2 = 4, RIGHT3 = 5;
parameter [3:0] LEFT1 = 6, LEFT2 = 7, LEFT3 = 8;
parameter [3:0] DOWN1 = 9, DOWN2 = 10, DOWN3 = 11;

parameter [0:40] map [0:40] = {
41'b11111111111111111111111111111111111111111,
41'b10000000000000000000000000000000000000001,
41'b10000000000000000000000000000000000000001,
41'b10000000000000000000000000000000000000001,
41'b10001111111111111110001111111111111110001,
41'b10001111111111111110001111111111111110001,
41'b10001111111111111110001111111111111110001,
41'b10001110000000000000000000000000001110001,
41'b10001110000000000000000000000000001110001,
41'b10001110000000000000000000000000001110001,
41'b10001110001111111111111111111110001110001,
41'b10001110001111111111111111111110001110001,
41'b10001110001111111111111111111110001110001,
41'b10001110000000000000000000000000001110001,
41'b10001110000000000000000000000000001110001,
41'b10001110000000000000000000000000001110001,
41'b10001110001111111111111111111111111110001,
41'b10001110001111111111111111111111111110001,
41'b10001110001111111111111111111111111110001,
41'b10001110000000000000000000000000000000000,
41'b10001110000000000000000000000000000000000,
41'b10001110000000000000000000000000000000000,
41'b10001110001111111111111111111111111110001,
41'b10001110001111111111111111111111111110001,
41'b10001110001111111111111111111111111110001,
41'b10001110001110000000000000000000001110001,
41'b10001110001110000000000000000000001110001,
41'b10001110001110000000000000000000001110001,
41'b10001110001110001110001110001110001110001,
41'b10001110001110001110001110001110001110001,
41'b10001110001110001110001110001110001110001,
41'b10000000000000001110001110001110001110001,
41'b10000000000000001110001110001110001110001,
41'b10000000000000001110001110001110001110001,
41'b11111111111111111111111110001110001110001,
41'b11111111111111111111111110001110001110001,
41'b11111111111111111111111110001110001110001,
41'b10000000000000000000000000001110000000001,
41'b10000000000000000000000000001110000000001,
41'b10000000000000000000000000001110000000001,
41'b11111111111111111111111111111111111111111
};

always @(posedge clk_23 or posedge rst) begin
    if (rst) player_state <= RIGHT1;
    else begin
        case(state)
        STAGE1, STAGE2, STAGE3: begin
            if(key_down[last_change]) begin
                case (key_num)
                4: player_state <= (player_state == UP2) ? UP3 : UP2;
                5: player_state <= (player_state == LEFT2) ? LEFT3 : LEFT2;
                6: player_state <= (player_state == DOWN2) ? DOWN3 : DOWN2;
                7: player_state <= (player_state == RIGHT2) ? RIGHT3 : RIGHT2;
                default: player_state <= player_state;
                endcase
            end else player_state <= player_state / 3 * 3;
        end
        default: player_state <= RIGHT1;
        endcase
    end
end

always @(posedge clk_23) begin
    player_x <= player_x;
    player_y <= player_y;
    case(state)
    STAGE1, STAGE2, STAGE3: begin
        if(key_down[last_change]) begin
            case (key_num)
            4: begin
                if(!map[(player_y -1 - 30)/5][(player_x - 60)/5] && !map[(player_y -1 - 30 +10)/5][(player_x - 60 +10)/5] && !map[(player_y -1 - 30+10)/5][(player_x - 60)/5] && !map[(player_y -1 - 30)/5][(player_x - 60 +10)/5])begin
                    player_y <= player_y - 1;
                end
            end
            5: begin
                if(!map[(player_y - 30)/5][(player_x -1 - 60)/5] && !map[(player_y - 30 +10)/5][(player_x -1 - 60 +10)/5] && !map[(player_y - 30+10)/5][(player_x -1 - 60)/5] && !map[(player_y - 30 )/5][(player_x -1 - 60 +10)/5])begin
                    player_x <= player_x - 1;
                end
            end
            6: begin
                if(!map[(player_y +1 - 30)/5][(player_x - 60)/5] && !map[(player_y +1 - 30 +10)/5][(player_x - 60 +10)/5] && !map[(player_y +1 - 30+10)/5][(player_x - 60)/5] && !map[(player_y +1 - 30 )/5][(player_x - 60 +10)/5])begin
                    player_y <= player_y + 1;
                end
            end
            7: begin
                if(!map[(player_y - 30)/5][(player_x +1 - 60)/5] && !map[(player_y - 30 +10)/5][(player_x +1 - 60 +10)/5] && !map[(player_y - 30+10)/5][(player_x +1 - 60)/5] && !map[(player_y - 30 )/5][(player_x +1 - 60 +10)/5])begin
                    player_x <= player_x + 1;
                end
            end
            endcase
        end
    end
    default: begin
        player_x <= 65;
        player_y <= 125;
    end
    endcase
end
//Boss position
reg [8:0] next_boss_x;
reg [8:0] next_boss_y;

parameter [0:337] shortest_dir[0:168]={
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10001111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000000000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000101000,
338'b10100011111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000000000000000000000000000000000001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000001000010101010101010100000101000,
338'b10101000111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000000000000000000000000000000000001111111111111000000000000010000000000000000001111111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010001111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000000000000000000000000000000000001111111111101000000000000010000000000010000001100111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010100011111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000000000000000000000000000000000001111111111101000000000000010000000000010000001000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101000111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000000000000000000000000000000000001111111111101000000000000010000000000010000001000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101010001111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111101010101000000000000000000000000000000000000001111111111001000000000000010000000000010000001000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101010100011111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111110101010101000000000000000000000000000000000000001111111101001000000000000010000000000010000001000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101010101000111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111010101010101000000000000000000000000000000000000001111110101001000000000000010000000000010000001000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101010101010001111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011101010101010101000000000000000000000000000000000000001111010101001000000000000010000000000010000001000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101010101010100011000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000010101010101010101000000000000000000000000000000000000001101010101001000000000000010000000000010000001000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101010101010101000000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000010101010101010101000000000000000000000000000000000000010101010101001000000000000010000000000010000001000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b01111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000111111111111110101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111110101000000000000000000000000000000000000001111111111111000000000000010000000000000000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101010101010101001000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000001010101010101010101000000000000000000000000000000000000010101010101001000000000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b01111111111111111111111111010000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000010000000000000000000000000111111111111111101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001100,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000001111111111111111000000000000000000000000000000000000111111111111110000000100000000000000000000000101000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000100011111111111111000000000000000000000000000000000000111111111111100000000000000000000000000000000001000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000101000111111111111000000000000000000000000000000000000111111111110100000000000000000000000000000000000000011111111111111111100010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000101010001111111111000000000000000000000000000000000000111111111010100000000000000000000000000000000000000011111111111111111000000000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000101000,
338'b10101010101001111111111111000000000000010000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111111101000000000000000000000000000000000000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000001000010101010101010100000101000,
338'b10101010101001111111111111000000000000010000000000000000101010101000111111000000000000000000000000000000000000111110101010100000000000000000000000000000000000000011111111111111101000000000000000000000000000000000000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000001000010101010101010100000101000,
338'b10101010101001111111111111000000000000010000000000000000101010101010001111000000000000000000000000000000000000111010101010100000000000000000000000000000000000000011111111111111101000000000000000000000000000000000000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000001000010101010101010100000101000,
338'b10101010101001111111111111000000000000010000000000000000101010101010100011000000000000000000000000000000000000101010101010100000000000000000000000000000000000000011111111111111101000000000000000000000000000000000000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000001000010101010101010100000101000,
338'b10101010101001111111111111000000000000010000000000000000101010101010101000000000000000000000000000000000000000101010101010100000000000000000000000000000000000000011111111111111101000000000000000000000000000000000000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000001000010101010101010100000101000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101010101010101001000000000000000000000000010000101010100011111111000000000000000000000000000000000000111111101010100000000000010000000000000000000000001010101010101010101000000000000000000000000000000000000010101010101001000001000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b01111111111111111111111111010000000000000000000000000100101010100011111111000000000000000000000000000000000001111111111010100000000000010000000000000000000000000111111111111111111000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000011111111111111111000000000000000000000000000000010000111111111111111100010100000000000000000000000101000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000101010101010101001000000000000000000000000000000000010101010101010100000000000000000000000000000000000000011111111111111111000000000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000101000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101010101010101001000000000000000000000000010000101010100011111111000100000000000000000000000000000001111111111010100000000000010000000000000000000000001010101010101010101000000000000000000000000000000100000010101010101001000001000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b01111111111111111111111111010000000000000000000000000100101010100011111111000001000100000000000000000000000001111111111110100000000000010000000000000000000000000111111111111111111100000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000011111111111111101000001000100000000000000010001010000111111111111111100010100000000000000000000000101000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000011111111111111001000001000100000000000000010001010010001111111111111100010100000000000000000000000101000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000011111111111101001000001000100000000000000010001010010100011111111111100010100000000000000000000000101000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000011111111110101001000001000100000000000000010001010010101000111111111100010100000000000000000000000101000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000011111111010101001000001000100000000000000010001010010101010001111111100010100000000000000000000000101000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000011111101010101001000000000100000000000000010000010010101010100011111100010100000000000000000000000101000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000011110101010101001000000000100000000000000010000000010101010101000111100000100000000000000000000000101000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000011010101010101001000000000100000000000000010000000010101010101010001100000000000000000000000000000001000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000000101010101010101001000000000100000000000000010000000010101010101010100000000000000000000000000000000000000011111111111111111100010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101010101010101001000000000000000000000000010000101010100011111111000100000100000000000000000001000001111111111110100000000000010000000000000000000000001010101010101010101000010000000000000000000000000100000010101010101001000001000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b01111111111111111111111111010000000000000000000000000100011010100011111111000001000100000000000000000000010001111111111111100000000000010000000000000000000000000111111111111111111111000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111111000000000000010000000000000100011111111111111101000101000100000000000000010001010001111111111111111100010100000000000000000000000101000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101010101010101001000000000000000000000000010000011010100011111111000100000100000000000000000001000001111111111111100000010000010000000000000000000001001010101010101010101000010000000000000000000000000100000010101010101001000001000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b01111111111111111111111111010000000000000000000000000100011110100011111111000001000100000000000000000000010001111111111111110000000100010000000000000000000100000111111111111111111111000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111101010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000011111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101001111111111001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101001000111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000101000,
338'b10101010101001111111101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101001010001111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000001000010101010101010100000101000,
338'b10101010101001111110101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101001010100011111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101001010101000111111111111010000000000000000000000000100000001111111111101000001000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101001101010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101001010101010001111111111010000000000000000000000000100000001111111111001000001000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101010101010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101001010101010100011111111010000000000000000000000000100000001111111101001000001000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101010101010101001000000000000000000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101001010101010101000111111010000000000000000000000000100000001111110101001000001000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101010101010101001000000000000000000000000010000011111110011111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101001010101010101010001111010000000000000000000000000100000001111010101001000001000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101010101010101001000000000000000000000000010000011111100011111111000100000100000000000000000001010001111111111111111100010100010000000000000000000101001010101010101010100011010000000000000000000000000100000001101010101001000001000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b10101010101010101010101001000000000000000000000000010000011110100011111111000100000100000000000000000001000001111111111111110000010100010000000000000000000101001010101010101010101000010000000000000000000000000100000010101010101001000001000000010000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b01111111111111111111111111010000000000000000000000000100011111100011111111000001000100000000000000000000010001111111111111111100010100010000000000000000000101000111111111111111111111000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01101010101001111111111101010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111111010000000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101010101010101001000000000000000000000000010000011110100011111111000100000100000000000000000001000001111111111111110000010100010000000000000000000101001010101010101010101001010000000000000000000000000100000010101010101001000001000000000000000000010000101000111100000000000100000000000000000000000001000010101010101010100000101000,
338'b01111111111111111111111111010000000000000000000000000100011111110011111101000001000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111111010001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01111010101001111111111101010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111111010001000000000000000000000100000001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001100,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01111111101001111111111101010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111101010001000000000000000000010100010000111111111111000101000100000000000000000001101010100000000000000000010000000000000000000000000110101010101010100000001111,
338'b01111111101001111111111001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111001010001000000000000000000010100010010001111111111000101000100000000000000000001101010100000000000000000010000000000000000000000000110101010101010100000001111,
338'b01111111101001111111101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111101001010001000000000000000000010100010010100011111111000101000100000000000000000001101010100000000000000000010000000000000000000000000110101010101010100000001111,
338'b01111111101001111110101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111110101001010001000000000000000000010100010010101000111111000101000100000000000000000001101010100000000000000000010000000000000000000000000110101010101010100000001111,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010001111000101000100000000000000000001101010100000000000000000010000000000000000000000000110101010101010100000001111,
338'b01111111101001101010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111101010101001010001000000000000000000010100010010101010100011000101000100000000000000000001101010100000000000000000010000000000000000000000000110101010101010100000001111,
338'b01111111101010101010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111110101010101001010001000000000000000000010100010010101010101000000101000100000000000000000001101010100000000000000000010000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101010101010101001000000000000000000000000010000011110100011111111000100000100000000000000000001000001111111111111110000010100010000000000000000000101001010101010101010101001010000000000000000000000010100000010101010101001000001000000000000000000010000101000110000000000000100000000000000000000000001000010101010101010100000101000,
338'b01111111111111111111111111010000000000000000000000000100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111111010001000000000000000000000100010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01111110101001111111111101010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111111010001000000000000000000000100010001111111111111000001000000010000000000000000101000111100000000000000000000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01111111101001111111111101010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111111010001000000000000000000000100010001111111111111000101000100000000000000000001101010100000000000000000010000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01111111101001111111101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111101001010001000000000000000000010100010010100111111111000101000100000000000000000001101010100000000000000000010000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000000000001101010100000000000000000010000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01111110101010101010101001010000000000000000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111010101010101001010001000000000000000000010100010010101010101001000101000100000000000000000001101010100000000000000000010000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101010101010101001000000000000000000000000010000011110100011111111000100000100000000000000000001000001111111111111110000010100010000000000000000000101001010101010101010101001010000000000000000000000010100000010101010101001000101000000000000000000010000101000100000000000000100000000000000000000000001000010101010101010100000101000,
338'b01111111111101111111111101010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111111010001000000000000000000000100010001111111111111000001000100010000000000000000001111111100000000000000000000000000000000000000000110101010101010100000001111,
338'b01111111111001111111111101010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111111010001000000000000000000000100010001111111111111000001000100010000000000000000100011111100000000000000000000000000000000000000000110101010101010100000001111,
338'b01111111101001111111111101010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111111010001000000000000000000000100010001111111111111000001000100010000000000000000101000111100000000000000000000000000000000000000000110101010101010100000001111,
338'b01111111101001111111111101010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111111010001000000000000000000000100010001111111111111000001000100010000000000000000101010001100000000000000010000000000000000000000000110101010101010100000001111,
338'b01111111101001111111111101010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111111111010001000000000000000000000100010001111111111111000001000100010000000000000001101010100000000000000000010000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01111111101001111111101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111111101001010001000000000000000000010100010010100111111111000101000100000001000000000001101010100000000000000000010000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000100000001101010100000000000000000010000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01111010101010101010101001010000000000000000000000010100011111110011111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111101010101010101001010001000000000000000000010100010010101010101001000101000100000000000000010001101010100000000000000000010000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101010101010101001000000000000000000000000010000011110100011111111000100000100000000000000000001000001111111111111110000010100010000000000000000000101001010101010101010101001010000000000000000000000010100000010101010101001000101000000000000000000010001101000100000000000000100000000000000000000000001001010101010101010100000101000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000100000001101010100000000001000000010000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b01101010101010101010101001010000000000000000000000010100011111100011111111000101000100000000000000000001010001111111111111111100010100010000000000000000000101000110101010101010101001010001000000000000000000010100010010101010101001000101000100000000000000010001101010100000000000000100010000000000000000000000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101010101010101001000000000000000000000000010000011110100011111111000100000100000000000000000001010001111111111111110000010100010000000000000000000101001010101010101010101001010000000000000000000000010100000010101010101001000101000000000000000000010001101010100000000000000100010000000000000000000001000010101010101010100000101000,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000100000001101010100000000001000000010000000000000000010000000100111111111111111100001111,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000100000001101010100000000001000000010000000000000000010000000110001111111111111100001111,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000100000001101010100000000001000000010000000000000000010000000110100011111111111100001111,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000100000001101010100000000001000000010000000000000000010000000110101000111111111100001111,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000100000001101010100000000001000000010000000000000000010000000110101010001111111100001111,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000100000001101010100000000001000000010000000000000000010000000110101010100011111100001111,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000100000001101010100000000001000000010000000000000000010000000110101010101000111100001111,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000100000001101010100000000001000000010000000000000000010000000110101010101010001100001111,
338'b01111111101001111010101001010000000000010000000000010100011111111111111101000101000100000000000000010001010001111111111111111100010100010000000000000000000101000111111111111010101001010001000000000000000000010100010010101010011111000101000100000000000100000001101010100000000001000000010000000000000000010000000010101010101010100000001111,
338'b00111111111111111111111111000000000000000000000000000000101010100011111111000000000000000000000000000000000000111111101010100000000000000000000000000000000000000011111111111010101000000001000000000000000000000000010001111111111111000000000100010000000000000000001111111100000000000000000000000000000000000000000010101010101010100000001000,
338'b10101010101010101010101001010000000000000000000000010100011110100011111111000101000100000000000000000001010001111111111111110000010100010000000000000000000101001010101010101010101001010001000000000000000000010100010010101010101001000101000100000000000000010001101010100000000000000100010000000000000000000001000110101010101010100000001111,
338'b10101010101010101010101001000000000000000000000000010100011110100011111111000101000100000000000000000001010001111111111111110000010100010000000000000000000101001010101010101010101001010000000000000000000000010100010010101010101001000101000100000000000000010001101010100000000000000100010000000000000000000001000110101010101010100000100011,
338'b10101010101010101010101001000000000000000000000000010000011110100011111111000101000100000000000000000001010001111111111111110000010100010000000000000000000101001010101010101010101001010000000000000000000000010100000010101010101001000101000100000000000000010001101010100000000000000100010000000000000000000001000110101010101010100000101000
};
//boss->player
wire [1:0] next_boss_dir;
reg [1:0] boss_dir;
wire [3:0] boss_x_maze ;
wire [3:0] boss_y_maze;
wire [3:0] player_x_maze ;
wire [3:0] player_y_maze ;
assign boss_x_maze = ((boss_x-60)/5-1)/3;
assign boss_y_maze = ((boss_y-30)/5-1)/3;
assign player_x_maze = ((player_x-60)/5-1)/3;
assign player_y_maze = ((player_y-30)/5-1)/3;
assign next_boss_dir = shortest_dir[(player_x_maze+player_y_maze*13)][(boss_x_maze+boss_y_maze*13)*2]*2+shortest_dir[(player_x_maze+player_y_maze*13)][(boss_x_maze+boss_y_maze*13)*2+1];
always @(posedge clk_23) begin
    if((boss_x-65)%15==2&&(boss_y-35)%15==2)begin
        boss_dir <= next_boss_dir;
    end
    else boss_dir<=boss_dir;
end
always @(posedge clk_23 or posedge rst) begin
    if (rst) boss_state <= RIGHT1;
    else begin
        case(state)
        STAGE3: begin
                case (boss_dir)
                0: boss_state <= (boss_state == UP2) ? UP3 : UP2;
                3: boss_state <= (boss_state == LEFT2) ? LEFT3 : LEFT2;
                1: boss_state <= (boss_state == DOWN2) ? DOWN3 : DOWN2;
                2: boss_state <= (boss_state == RIGHT2) ? RIGHT3 : RIGHT2;
                default: boss_state <= boss_state;
                endcase
        end
        default: boss_state <= RIGHT1;
        endcase
    end
end
always @(posedge clk_23 or posedge rst) begin
    if(rst)begin
        boss_x <=  247;
        boss_y <= 37;
    end
    else begin
        boss_x <=  boss_x;
        boss_y <= boss_y;
        
        case(state)
        STAGE3:begin
        case (boss_dir)
            0: begin
                if(!map[(boss_y -1 - 30)/5][(boss_x - 60)/5] && !map[(boss_y -1 - 30 +10)/5][(boss_x - 60 +10)/5])begin
                    boss_y <= boss_y - 1;
                end
            end
            3: begin
                if(!map[(boss_y - 30)/5][(boss_x -1 - 60)/5] && !map[(boss_y - 30 +10)/5][(boss_x -1 - 60 +10)/5])begin
                    boss_x <= boss_x - 1;
                end
            end
            1: begin
                if(!map[(boss_y +1 - 30)/5][(boss_x - 60)/5] && !map[(boss_y +1 - 30 +10)/5][(boss_x - 60 +10)/5])begin
                    boss_y <= boss_y + 1;
                end
            end
            2: begin
                if(!map[(boss_y - 30)/5][(boss_x +1 - 60)/5] && !map[(boss_y - 30 +10)/5][(boss_x +1 - 60 +10)/5])begin
                    boss_x <= boss_x + 1;
                end
            end
            endcase
        end
        endcase
    end
end

// Object Position

// Collide
// Key
always @(posedge clk_23) begin
    key_find <= key_find;
    case(state)
    STAGE1, STAGE3: begin
        case (key_find)
        0: begin
            if (player_x >= 55 && player_x < 85 && player_y >= 25 && player_y < 55)
                key_find <= key_find + 1;
        end
        1: begin
            if (player_x >= 220 && player_x < 250 && player_y >= 25 && player_y < 55)
                key_find <= key_find + 1;
        end
        2: begin
            if (player_x >= 220 && player_x < 250 && player_y >= 195 && player_y < 255)
                key_find <= key_find + 1;
        end
        endcase
    end
    STAGE2: begin
        if (!isDark) begin
            case (key_find)
            0: begin
                if (player_x >= 55 && player_x < 85 && player_y >= 25 && player_y < 55)
                    key_find <= key_find + 1;
            end
            1: begin
                if (player_x >= 220 && player_x < 250 && player_y >= 25 && player_y < 55)
                    key_find <= key_find + 1;
            end
            2: begin
                if (player_x >= 220 && player_x < 250 && player_y >= 195 && player_y < 255)
                    key_find <= key_find + 1;
            end
            endcase
        end
    end
    default: key_find <= 0;
    endcase
end
// Pass
always @(posedge clk_23) begin
    if (key_find == 3 && player_x >= 250 && player_x < 280 && player_y >= 110 && player_y < 140)
        pass <= 1;
    else pass <= 0;
end
// Light
always @(posedge clk_23) begin
    isDark <= isDark;
    case(state)
    STAGE2: begin
        if (player_x >= 170 && player_x < 200 && player_y >= 125 && player_y < 150)
            isDark <= 0;
    end
    default: isDark <= 1;
    endcase
end
endmodule

