// wall
`define wall_h = 0;
`define wall_v = 20;

`define rec_h = 10;
`define rec_v = 10; 
module draw_interface(
    input [3:0] state;
    input [9:0] h_cnt;
    input [9:0] v_cnt;
    input [1:0] key_find;
    output [16:0] pixel_addr;
)
parameter [3:0] TITLE = 0, STAFF = 1;
parameter [3:0] STAGE1 = 2, SUCCESS1 = 3;
parameter [3:0] STAGE2 = 4, SUCCESS2 = 5;
parameter [3:0] STAGE3 = 6, SUCCESS3 = 7, FAIL = 8;

parameter [39:0] map [39:0] = {
    40'b111111111111111111111111111111111111111,
    40'b100000000000000000010000000000000000001,
    40'b100000000000000000010000000000000000001,
    40'b100000000000000000010000000000000000001,
    40'b100000000000000000010000000000000000001,
    40'b100001111111111000011111111111111100001,
    40'b100001000000000000000000000000000100001,
    40'b100001000000000000000000000000000100001,
    40'b100001000000000000000000000000000100001,
    40'b100001000000000000000000000000000100001,
    40'b100001000011111111111111111110000100001,
    40'b100001000000000000000000000000000100001,
    40'b100001000000000000000000000000000100001,
    40'b100001000000000000000000000000000100001,
    40'b100001000000000000000000000000000100001,
    40'b100001000011111111111111111111111100001,
    40'b100001000000000000000000000000000000000,
    40'b100001000000000000000000000000000000000,
    40'b000001000000000000000000000000000000000,
    40'b000001000000000000000000000000000000000,
    40'b000001000011111111111111111111111100001,
    40'b000001000010000000000000000000000100001,
    40'b100001000010000000000000000000000100001,
    40'b100001000010000000000000000000000100001,
    40'b100001000010000000000000000000000100001,
    40'b100001000010000100001100001000000100001,
    40'b100001000010000100001100001000000000001,
    40'b100001000010000100001100001000000000001,
    40'b100001000010000100001100001000000000001,
    40'b100000000000000100001100001000000000001,
    40'b100000000000000100001100001000011100001,
    40'b100000000000000100001100001000011100001,
    40'b100000000000000100001100001000011100001,
    40'b111111111111111111111100001000011100001,
    40'b111111111111111111111100001000011100001,
    40'b100000000000000000000000001000000000001,
    40'b100000000000000000000000001000000000001,
    40'b100000000000000000000000001000000000001,
    40'b100000000000000000000000001000000000001,
    40'b111111111111111111111111111111111111111
};
wire [8:0] x,y;
assign x = (h_cnt<<1);
assign y = (v_cnt<<1);
always@(*)begin
    case(state)
    STAGE1:begin
        if(map[x/5][y/5])begin
            pixel_addr = (x%5+(y%5+120)*320)%76800;
        end
    end
    endcase
end
endmodule
//200*200->40*40 player20*20->4*4
/*

111111111111111111111111111111111111111
100000000000000000010000000000000000001
100000000000000000010000000000000000001
100000000000000000010000000000000000001
100000000000000000010000000000000000001
100001111111111000011111111111111100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000011111111111111111110000100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000000000000000000000000000100001
100001000011111111111111111111111100001
100001000000000000000000000000000000000
100001000000000000000000000000000000000
000001000000000000000000000000000000000
000001000000000000000000000000000000000
000001000011111111111111111111111100001
000001000010000000000000000000000100001
100001000010000000000000000000000100001
100001000010000000000000000000000100001
100001000010000000000000000000000100001
100001000010000100001100001000000100001
100001000010000100001100001000000000001
100001000010000100001100001000000000001
100001000010000100001100001000000000001
100000000000000100001100001000000000001
100000000000000100001100001000011100001
100000000000000100001100001000011100001
100000000000000100001100001000011100001
111111111111111111111100001000011100001
111111111111111111111100001000011100001
100000000000000000000000001000000000001
100000000000000000000000001000000000001
100000000000000000000000001000000000001
100000000000000000000000001000000000001
111111111111111111111111111111111111111
*/